// (c) Technion IIT, Department of Electrical Engineering 2022 
// Updated by Mor Dahan - January 2022


module time_place_word 
	(
	output	[10:0] xPos_1,
	output	[10:0] yPos_1
	
	); 
	
assign xPos = 64;
assign yPos = 32;

endmodule 