// System-Verilog 'written by Alex Grinshpun May 2018
// New bitmap dudy February 2021
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	mineMatrixBitMap_v2	(		
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic mine_Collision,

					output	logic	minedrawingRequest, //output that a mine would be dispalyed
					output	logic	[7:0] RGBout, 
					output   logic mine_exploded //block_broken
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */
 logic [3:0] Block_To_Break_Y;
 logic [4:0] Block_To_Break_X;

// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 



logic [0:14] [0:19] [3:0]  MazeBiMapMask= 
{{4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h01, 4'h01, 4'h01, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h01, 4'h01, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
 {4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01}};

 
 
logic [0:31] [0:31] [7:0]  object_colors  ={
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h24,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'h00,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'h00,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'h00,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'h00,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'h00,8'hfe,8'hb5,8'hb1,8'hb1,8'hb1,8'hfe,8'hfa,8'hfe,8'hfe,8'hd5,8'hfe,8'hb1,8'hb1,8'hb1,8'hfa,8'hfe,8'h00,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'h00,8'h00,8'h00,8'h00,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'h00,8'h00,8'h00,8'h00,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hfc,8'hfc,8'hfc,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'h00,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'hfc,8'hfc,8'hfc,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hfc,8'hfc,8'hfc,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'hff,8'h00,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'hfc,8'hfc,8'hfc,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'h00,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'hfe,8'h00,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'h00,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'h00,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'h00,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'h00,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'ha4,8'hec,8'hff,8'hec,8'hec,8'hec,8'h00,8'hec,8'hff,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'h00,8'hec,8'hec,8'hec,8'hec,8'hec,8'h00,8'hec,8'hec,8'hec,8'hec,8'he0,8'h00,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hff,8'hff,8'hff}};




// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
		MazeBiMapMask <= 
		{{4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h05, 4'h05, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
		 {4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h01, 4'h01, 4'h01, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h04, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h03, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h03, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h06, 4'h06, 4'h03, 4'h01, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01},
		 {4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01, 4'h01}};
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
		   (MazeBiMapMask[offsetY[8:5]][offsetX[9:5]] == 4'h01 )) // take bits 5,6,7,8,9,10 from address to select  position in the maze    
						RGBout <= object_colors[4'h00][offsetY[4:0]][offsetX[4:0]] ;
						
		
		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
		   (MazeBiMapMask[offsetY[8:5] ][offsetX[9:5]] == 4'h01 ) & (mine_Collision)) // take bits 5,6,7,8,9,10 from address to select  position in the maze    
						MazeBiMapMask[offsetY[8:5] ][offsetX[9:5]] <= 4'h00 ;
						mine_exploded=1'b1;
						
		end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 

assign minedrawingRequest = ((RGBout != TRANSPARENT_ENCODING) && (MazeBiMapMask[offsetY[8:5]][offsetX[9:5]] == 4'h01)) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap


endmodule


