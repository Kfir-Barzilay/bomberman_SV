// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen Apr  	0	3  
// (c) Technion IIT, Department of Electrical Engineering 	0	3 



module	HartsMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic [7:0] random_hart,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  	0 * 15 squares of 3	*3	  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares 
// this is the bitmap  of the maze , if there is a specific value  the  whole 3	*3	 rectange will be drawn on the screen
// there are  16 options of differents kinds of 32*32 squares 
// all numbers here are hard coded to simplify the  understanding 



logic [0:12] [0:17] [3:0]  MazeBiMapMask= 
{{4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00},
 {4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00},
 {4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00},
 {4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00},
 {4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00},
 {4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00, 4'h01, 4'h00},
 {4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h00, 4'h01, 4'h00}};


 logic [0:2] [0:31] [0:31] [7:0]  object_colors  = {
  {{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d}}
,  {
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h91,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h91,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h91,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'hb6,8'h00,8'h91,8'h91},
	{8'h91,8'hb6,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'hb6,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h91,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h91,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h91,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'hb6,8'h00,8'h91,8'h91},
	{8'h91,8'hb6,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'hb6,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h91,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h91,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h91,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'hb6,8'h00,8'h91,8'h91},
	{8'h91,8'hb6,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'hb6,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h91,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h91,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h91,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'hb6,8'h00,8'h91,8'h91},
	{8'h91,8'hb6,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'hb6,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d}}

 
, {
	{8'h8d,8'h65,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h8d,8'h00,8'h8d,8'h64,8'h6d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h8d,8'h00,8'h8d,8'h65,8'h8d,8'h8d,8'h00,8'h8d,8'h65,8'h8d,8'h8d,8'h00,8'h8d,8'h64},
	{8'h8d,8'h8d,8'h8d,8'h8d,8'h00,8'h6d,8'h8d,8'h8d,8'h6d,8'h00,8'h8d,8'h8d,8'h8d,8'h6d,8'h00,8'h8d,8'h8d,8'h8d,8'h8d,8'h00,8'h8d,8'h8d,8'h6d,8'h8d,8'h00,8'h8d,8'h8d,8'h8d,8'h8d,8'h00,8'h8d,8'h8d},
	{8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'hb1,8'h64,8'hb1,8'h91,8'h00,8'hb1,8'h64,8'hb1,8'hb1,8'h00,8'hb1,8'h64,8'hb1,8'h91,8'h00,8'hb1,8'h64,8'hb1,8'h91,8'h00,8'hb1,8'h65,8'h91,8'h91,8'h00,8'h91,8'h64,8'hb1,8'h91,8'h00,8'hb2,8'h65},
	{8'hb1,8'hb2,8'hb1,8'h91,8'h00,8'h91,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'hb1,8'h91,8'h91,8'h00,8'hb1,8'h91,8'hb2,8'h91,8'h00,8'h91,8'h91,8'h95,8'h91,8'h00,8'hb6,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91},
	{8'hb1,8'h91,8'hb1,8'h91,8'h00,8'h91,8'hb1,8'hb1,8'h91,8'h00,8'hb2,8'hb1,8'h91,8'h91,8'h00,8'hb1,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'hb1},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h8d,8'h65,8'h6d,8'h6d,8'h00,8'h6d,8'h65,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h8d,8'h00,8'h8d,8'h65,8'h6d,8'h6d,8'h00,8'h6d,8'h64,8'h8d,8'h8d,8'h00,8'h8d,8'h64},
	{8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h8d,8'h8d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h8d,8'h00,8'h6d,8'h6d,8'h6d,8'h8d,8'h00,8'h6d,8'h6d,8'h8d,8'h6d,8'h00,8'h8d,8'h6d},
	{8'h8d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h8d,8'h8d,8'h6d,8'h00,8'h6d,8'h8d,8'h71,8'h6d,8'h00,8'h6d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h8d,8'h6d,8'h6d,8'h8d,8'h00,8'h6d,8'h6d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'hb1,8'h64,8'h91,8'h96,8'h00,8'h91,8'h64,8'hb1,8'h91,8'h00,8'hb2,8'h64,8'hb1,8'h91,8'h00,8'hb1,8'h64,8'hb1,8'hb1,8'h00,8'hb1,8'h65,8'h91,8'h91,8'h00,8'h91,8'h6d,8'hb1,8'h91,8'h00,8'hb1,8'h64},
	{8'hb1,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'h91,8'hb1,8'h91,8'h00,8'hb1,8'h91,8'h91,8'h91,8'h00,8'h91,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'hb1,8'h91,8'h91,8'h00,8'h91,8'hb2},
	{8'hb1,8'hb1,8'hb1,8'h91,8'h00,8'hb1,8'hb1,8'hb1,8'hb1,8'h00,8'hb1,8'hb1,8'h91,8'h91,8'h00,8'h91,8'hb1,8'hb1,8'h91,8'h00,8'hb1,8'hb1,8'h91,8'h91,8'h00,8'h91,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h6d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64},
	{8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h8d,8'h8d,8'h6d,8'h00,8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h8d,8'h6d,8'h00,8'h8d,8'h8d},
	{8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h8d,8'h6d,8'h6d,8'h00,8'h8d,8'h8d,8'h91,8'h6d,8'h00,8'h6d,8'h8d,8'h6d,8'h6d,8'h00,8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h8d,8'h8d,8'h6d,8'h00,8'h6d,8'h8d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'hb1,8'h64,8'h91,8'hb6,8'h00,8'hb1,8'h64,8'hb1,8'h91,8'h00,8'hb2,8'h64,8'hb1,8'h91,8'h00,8'hb1,8'h64,8'hb1,8'h91,8'h00,8'hb1,8'h65,8'h91,8'h91,8'h00,8'h91,8'h65,8'hb1,8'h91,8'h00,8'hb1,8'h64},
	{8'hb1,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'h91,8'hb1,8'h91,8'h00,8'h91,8'h91,8'hb1,8'h91,8'h00,8'h91,8'h91,8'hb1,8'h91,8'h00,8'h91,8'h91,8'h91,8'hb1,8'h00,8'h91,8'hb1,8'h91,8'h91,8'h00,8'h91,8'hb2},
	{8'hb1,8'h91,8'h91,8'hb1,8'h00,8'hb1,8'hb1,8'hb1,8'hb1,8'h00,8'hb1,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'hb1,8'h91,8'h91,8'h00,8'h91,8'hb1,8'hb1,8'hb1,8'h00,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h6d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64},
	{8'h6d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h6d,8'h6d,8'h8d,8'h6d,8'h00,8'h8d,8'h8d},
	{8'h8d,8'h6d,8'h6d,8'h6d,8'h00,8'h6d,8'h91,8'h6d,8'h6d,8'h00,8'h6d,8'h8d,8'h91,8'h6d,8'h00,8'h6d,8'h8d,8'h6d,8'h6d,8'h00,8'h8d,8'h8d,8'h6d,8'h6d,8'h00,8'h8d,8'h8d,8'h8d,8'h6d,8'h00,8'h6d,8'h8d},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'hb1,8'h64,8'h91,8'h96,8'h00,8'hb1,8'h64,8'hb1,8'h91,8'h00,8'hb2,8'h64,8'hb1,8'h91,8'h00,8'hb1,8'h64,8'hb1,8'hb1,8'h00,8'hb1,8'h65,8'h91,8'h91,8'h00,8'h91,8'h6d,8'hb1,8'h91,8'h00,8'hb1,8'h64},
	{8'hb1,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'h91,8'hb1,8'h91,8'h00,8'hb1,8'h91,8'hb1,8'h91,8'h00,8'h91,8'h91,8'hb1,8'hb1,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'h91,8'h00,8'h91,8'hb2},
	{8'hb1,8'h91,8'h91,8'hb1,8'h00,8'hb1,8'hb1,8'hb1,8'hb1,8'h00,8'hb1,8'hb1,8'hb1,8'h91,8'h00,8'h91,8'h91,8'hb1,8'h91,8'h00,8'h91,8'hb1,8'h91,8'h91,8'h00,8'h91,8'h91,8'h91,8'hb1,8'h00,8'h91,8'h91},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h6d,8'h00,8'h8d,8'h64,8'h8d,8'h8d,8'h00,8'h8d,8'h64,8'h8d,8'h8d,8'h00,8'h8d,8'h64,8'h8d,8'h8d,8'h00,8'h8d,8'h64}}

 };
 

// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
		   (MazeBiMapMask[offsetY[8:5] ][offsetX[8:5]] == 4'h01 )) // take bits 5,6,7,8,9,10 from address to select  position in the maze    
						RGBout <= object_colors[2'b10][offsetY[4:0]][offsetX[4:0]] ; 
		end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule

